`timescale 1ns / 1ps

`include "incl.vh"

//
// Provide w for compression loop instants.
//
module w_shift (
    input clk,
    input [511:0] chunk,
    output [32*64-1:0] out_w
);  
    //
    // w[0..15]
    //
    genvar k;
    wire [32*64-1:0] w;

    generate
        for (k=0; k<16; k=k+1) begin
            w_0_15 #(
                .DELAY_OUT_W(k*4)
            ) w_0_15_inst(
            	.clk(clk),
                .chunk(chunk[32*k+:32]),
                .out_w(w[32*k+:32]),
                .out_w_delayed(out_w[32*k+:32])
            );
        end
    endgenerate

    //
    // w[16..63], generated by gen_w_inst
    //
    w_16_63 #(  // w16, inputs should be aligned
        .DELAY_DIST_16(0),  // w0, delay 0 cycles
        .DELAY_DIST_15(0),  // w1, delay 0 cycles
        .DELAY_DIST_7(0),  // w9, delay 0 cycles
        .DELAY_DIST_2(0),  // w14, delay 0 cycles
        .DELAY_OUT_W(61)
    ) w_16_inst( 
        .clk(clk),
        .dist_16(w[31:0]),  // w0
        .dist_15(w[63:32]),  // w1
        .dist_7(w[319:288]),  // w9
        .dist_2(w[479:448]),  // w14
        .out_w(w[543:512]),
        .out_w_delayed(out_w[543:512])
    );

    w_16_63 #(  // w17, inputs should be aligned
        .DELAY_DIST_16(0),  // w1, delay 0 cycles
        .DELAY_DIST_15(0),  // w2, delay 0 cycles
        .DELAY_DIST_7(0),  // w10, delay 0 cycles
        .DELAY_DIST_2(0),  // w15, delay 0 cycles
        .DELAY_OUT_W(65)
    ) w_17_inst( 
        .clk(clk),
        .dist_16(w[63:32]),  // w1
        .dist_15(w[95:64]),  // w2
        .dist_7(w[351:320]),  // w10
        .dist_2(w[511:480]),  // w15
        .out_w(w[575:544]),
        .out_w_delayed(out_w[575:544])
    );

    w_16_63 #(  // w18, inputs should be aligned
        .DELAY_DIST_16(3),  // w2, delay 3 cycles
        .DELAY_DIST_15(3),  // w3, delay 3 cycles
        .DELAY_DIST_7(3),  // w11, delay 3 cycles
        .DELAY_DIST_2(0),  // w16, delay 0 cycles
        .DELAY_OUT_W(66)
    ) w_18_inst( 
        .clk(clk),
        .dist_16(w[95:64]),  // w2
        .dist_15(w[127:96]),  // w3
        .dist_7(w[383:352]),  // w11
        .dist_2(w[543:512]),  // w16
        .out_w(w[607:576]),
        .out_w_delayed(out_w[607:576])
    );

    w_16_63 #(  // w19, inputs should be aligned
        .DELAY_DIST_16(3),  // w3, delay 3 cycles
        .DELAY_DIST_15(3),  // w4, delay 3 cycles
        .DELAY_DIST_7(3),  // w12, delay 3 cycles
        .DELAY_DIST_2(0),  // w17, delay 0 cycles
        .DELAY_OUT_W(70)
    ) w_19_inst( 
        .clk(clk),
        .dist_16(w[127:96]),  // w3
        .dist_15(w[159:128]),  // w4
        .dist_7(w[415:384]),  // w12
        .dist_2(w[575:544]),  // w17
        .out_w(w[639:608]),
        .out_w_delayed(out_w[639:608])
    );

    w_16_63 #(  // w20, inputs should be aligned
        .DELAY_DIST_16(6),  // w4, delay 6 cycles
        .DELAY_DIST_15(6),  // w5, delay 6 cycles
        .DELAY_DIST_7(6),  // w13, delay 6 cycles
        .DELAY_DIST_2(0),  // w18, delay 0 cycles
        .DELAY_OUT_W(71)
    ) w_20_inst( 
        .clk(clk),
        .dist_16(w[159:128]),  // w4
        .dist_15(w[191:160]),  // w5
        .dist_7(w[447:416]),  // w13
        .dist_2(w[607:576]),  // w18
        .out_w(w[671:640]),
        .out_w_delayed(out_w[671:640])
    );

    w_16_63 #(  // w21, inputs should be aligned
        .DELAY_DIST_16(6),  // w5, delay 6 cycles
        .DELAY_DIST_15(6),  // w6, delay 6 cycles
        .DELAY_DIST_7(6),  // w14, delay 6 cycles
        .DELAY_DIST_2(0),  // w19, delay 0 cycles
        .DELAY_OUT_W(75)
    ) w_21_inst( 
        .clk(clk),
        .dist_16(w[191:160]),  // w5
        .dist_15(w[223:192]),  // w6
        .dist_7(w[479:448]),  // w14
        .dist_2(w[639:608]),  // w19
        .out_w(w[703:672]),
        .out_w_delayed(out_w[703:672])
    );

    w_16_63 #(  // w22, inputs should be aligned
        .DELAY_DIST_16(9),  // w6, delay 9 cycles
        .DELAY_DIST_15(9),  // w7, delay 9 cycles
        .DELAY_DIST_7(9),  // w15, delay 9 cycles
        .DELAY_DIST_2(0),  // w20, delay 0 cycles
        .DELAY_OUT_W(76)
    ) w_22_inst( 
        .clk(clk),
        .dist_16(w[223:192]),  // w6
        .dist_15(w[255:224]),  // w7
        .dist_7(w[511:480]),  // w15
        .dist_2(w[671:640]),  // w20
        .out_w(w[735:704]),
        .out_w_delayed(out_w[735:704])
    );

    w_16_63 #(  // w23, inputs should be aligned
        .DELAY_DIST_16(9),  // w7, delay 9 cycles
        .DELAY_DIST_15(9),  // w8, delay 9 cycles
        .DELAY_DIST_7(6),  // w16, delay 6 cycles
        .DELAY_DIST_2(0),  // w21, delay 0 cycles
        .DELAY_OUT_W(80)
    ) w_23_inst( 
        .clk(clk),
        .dist_16(w[255:224]),  // w7
        .dist_15(w[287:256]),  // w8
        .dist_7(w[543:512]),  // w16
        .dist_2(w[703:672]),  // w21
        .out_w(w[767:736]),
        .out_w_delayed(out_w[767:736])
    );

    w_16_63 #(  // w24, inputs should be aligned
        .DELAY_DIST_16(12),  // w8, delay 12 cycles
        .DELAY_DIST_15(12),  // w9, delay 12 cycles
        .DELAY_DIST_7(9),  // w17, delay 9 cycles
        .DELAY_DIST_2(0),  // w22, delay 0 cycles
        .DELAY_OUT_W(81)
    ) w_24_inst( 
        .clk(clk),
        .dist_16(w[287:256]),  // w8
        .dist_15(w[319:288]),  // w9
        .dist_7(w[575:544]),  // w17
        .dist_2(w[735:704]),  // w22
        .out_w(w[799:768]),
        .out_w_delayed(out_w[799:768])
    );

    w_16_63 #(  // w25, inputs should be aligned
        .DELAY_DIST_16(12),  // w9, delay 12 cycles
        .DELAY_DIST_15(12),  // w10, delay 12 cycles
        .DELAY_DIST_7(6),  // w18, delay 6 cycles
        .DELAY_DIST_2(0),  // w23, delay 0 cycles
        .DELAY_OUT_W(85)
    ) w_25_inst( 
        .clk(clk),
        .dist_16(w[319:288]),  // w9
        .dist_15(w[351:320]),  // w10
        .dist_7(w[607:576]),  // w18
        .dist_2(w[767:736]),  // w23
        .out_w(w[831:800]),
        .out_w_delayed(out_w[831:800])
    );

    w_16_63 #(  // w26, inputs should be aligned
        .DELAY_DIST_16(15),  // w10, delay 15 cycles
        .DELAY_DIST_15(15),  // w11, delay 15 cycles
        .DELAY_DIST_7(9),  // w19, delay 9 cycles
        .DELAY_DIST_2(0),  // w24, delay 0 cycles
        .DELAY_OUT_W(86)
    ) w_26_inst( 
        .clk(clk),
        .dist_16(w[351:320]),  // w10
        .dist_15(w[383:352]),  // w11
        .dist_7(w[639:608]),  // w19
        .dist_2(w[799:768]),  // w24
        .out_w(w[863:832]),
        .out_w_delayed(out_w[863:832])
    );

    w_16_63 #(  // w27, inputs should be aligned
        .DELAY_DIST_16(15),  // w11, delay 15 cycles
        .DELAY_DIST_15(15),  // w12, delay 15 cycles
        .DELAY_DIST_7(6),  // w20, delay 6 cycles
        .DELAY_DIST_2(0),  // w25, delay 0 cycles
        .DELAY_OUT_W(90)
    ) w_27_inst( 
        .clk(clk),
        .dist_16(w[383:352]),  // w11
        .dist_15(w[415:384]),  // w12
        .dist_7(w[671:640]),  // w20
        .dist_2(w[831:800]),  // w25
        .out_w(w[895:864]),
        .out_w_delayed(out_w[895:864])
    );

    w_16_63 #(  // w28, inputs should be aligned
        .DELAY_DIST_16(18),  // w12, delay 18 cycles
        .DELAY_DIST_15(18),  // w13, delay 18 cycles
        .DELAY_DIST_7(9),  // w21, delay 9 cycles
        .DELAY_DIST_2(0),  // w26, delay 0 cycles
        .DELAY_OUT_W(91)
    ) w_28_inst( 
        .clk(clk),
        .dist_16(w[415:384]),  // w12
        .dist_15(w[447:416]),  // w13
        .dist_7(w[703:672]),  // w21
        .dist_2(w[863:832]),  // w26
        .out_w(w[927:896]),
        .out_w_delayed(out_w[927:896])
    );

    w_16_63 #(  // w29, inputs should be aligned
        .DELAY_DIST_16(18),  // w13, delay 18 cycles
        .DELAY_DIST_15(18),  // w14, delay 18 cycles
        .DELAY_DIST_7(6),  // w22, delay 6 cycles
        .DELAY_DIST_2(0),  // w27, delay 0 cycles
        .DELAY_OUT_W(95)
    ) w_29_inst( 
        .clk(clk),
        .dist_16(w[447:416]),  // w13
        .dist_15(w[479:448]),  // w14
        .dist_7(w[735:704]),  // w22
        .dist_2(w[895:864]),  // w27
        .out_w(w[959:928]),
        .out_w_delayed(out_w[959:928])
    );

    w_16_63 #(  // w30, inputs should be aligned
        .DELAY_DIST_16(21),  // w14, delay 21 cycles
        .DELAY_DIST_15(21),  // w15, delay 21 cycles
        .DELAY_DIST_7(9),  // w23, delay 9 cycles
        .DELAY_DIST_2(0),  // w28, delay 0 cycles
        .DELAY_OUT_W(96)
    ) w_30_inst( 
        .clk(clk),
        .dist_16(w[479:448]),  // w14
        .dist_15(w[511:480]),  // w15
        .dist_7(w[767:736]),  // w23
        .dist_2(w[927:896]),  // w28
        .out_w(w[991:960]),
        .out_w_delayed(out_w[991:960])
    );

    w_16_63 #(  // w31, inputs should be aligned
        .DELAY_DIST_16(21),  // w15, delay 21 cycles
        .DELAY_DIST_15(18),  // w16, delay 18 cycles
        .DELAY_DIST_7(6),  // w24, delay 6 cycles
        .DELAY_DIST_2(0),  // w29, delay 0 cycles
        .DELAY_OUT_W(100)
    ) w_31_inst( 
        .clk(clk),
        .dist_16(w[511:480]),  // w15
        .dist_15(w[543:512]),  // w16
        .dist_7(w[799:768]),  // w24
        .dist_2(w[959:928]),  // w29
        .out_w(w[1023:992]),
        .out_w_delayed(out_w[1023:992])
    );

    w_16_63 #(  // w32, inputs should be aligned
        .DELAY_DIST_16(21),  // w16, delay 21 cycles
        .DELAY_DIST_15(21),  // w17, delay 21 cycles
        .DELAY_DIST_7(9),  // w25, delay 9 cycles
        .DELAY_DIST_2(0),  // w30, delay 0 cycles
        .DELAY_OUT_W(101)
    ) w_32_inst( 
        .clk(clk),
        .dist_16(w[543:512]),  // w16
        .dist_15(w[575:544]),  // w17
        .dist_7(w[831:800]),  // w25
        .dist_2(w[991:960]),  // w30
        .out_w(w[1055:1024]),
        .out_w_delayed(out_w[1055:1024])
    );

    w_16_63 #(  // w33, inputs should be aligned
        .DELAY_DIST_16(21),  // w17, delay 21 cycles
        .DELAY_DIST_15(18),  // w18, delay 18 cycles
        .DELAY_DIST_7(6),  // w26, delay 6 cycles
        .DELAY_DIST_2(0),  // w31, delay 0 cycles
        .DELAY_OUT_W(105)
    ) w_33_inst( 
        .clk(clk),
        .dist_16(w[575:544]),  // w17
        .dist_15(w[607:576]),  // w18
        .dist_7(w[863:832]),  // w26
        .dist_2(w[1023:992]),  // w31
        .out_w(w[1087:1056]),
        .out_w_delayed(out_w[1087:1056])
    );

    w_16_63 #(  // w34, inputs should be aligned
        .DELAY_DIST_16(21),  // w18, delay 21 cycles
        .DELAY_DIST_15(21),  // w19, delay 21 cycles
        .DELAY_DIST_7(9),  // w27, delay 9 cycles
        .DELAY_DIST_2(0),  // w32, delay 0 cycles
        .DELAY_OUT_W(106)
    ) w_34_inst( 
        .clk(clk),
        .dist_16(w[607:576]),  // w18
        .dist_15(w[639:608]),  // w19
        .dist_7(w[895:864]),  // w27
        .dist_2(w[1055:1024]),  // w32
        .out_w(w[1119:1088]),
        .out_w_delayed(out_w[1119:1088])
    );

    w_16_63 #(  // w35, inputs should be aligned
        .DELAY_DIST_16(21),  // w19, delay 21 cycles
        .DELAY_DIST_15(18),  // w20, delay 18 cycles
        .DELAY_DIST_7(6),  // w28, delay 6 cycles
        .DELAY_DIST_2(0),  // w33, delay 0 cycles
        .DELAY_OUT_W(110)
    ) w_35_inst( 
        .clk(clk),
        .dist_16(w[639:608]),  // w19
        .dist_15(w[671:640]),  // w20
        .dist_7(w[927:896]),  // w28
        .dist_2(w[1087:1056]),  // w33
        .out_w(w[1151:1120]),
        .out_w_delayed(out_w[1151:1120])
    );

    w_16_63 #(  // w36, inputs should be aligned
        .DELAY_DIST_16(21),  // w20, delay 21 cycles
        .DELAY_DIST_15(21),  // w21, delay 21 cycles
        .DELAY_DIST_7(9),  // w29, delay 9 cycles
        .DELAY_DIST_2(0),  // w34, delay 0 cycles
        .DELAY_OUT_W(111)
    ) w_36_inst( 
        .clk(clk),
        .dist_16(w[671:640]),  // w20
        .dist_15(w[703:672]),  // w21
        .dist_7(w[959:928]),  // w29
        .dist_2(w[1119:1088]),  // w34
        .out_w(w[1183:1152]),
        .out_w_delayed(out_w[1183:1152])
    );

    w_16_63 #(  // w37, inputs should be aligned
        .DELAY_DIST_16(21),  // w21, delay 21 cycles
        .DELAY_DIST_15(18),  // w22, delay 18 cycles
        .DELAY_DIST_7(6),  // w30, delay 6 cycles
        .DELAY_DIST_2(0),  // w35, delay 0 cycles
        .DELAY_OUT_W(115)
    ) w_37_inst( 
        .clk(clk),
        .dist_16(w[703:672]),  // w21
        .dist_15(w[735:704]),  // w22
        .dist_7(w[991:960]),  // w30
        .dist_2(w[1151:1120]),  // w35
        .out_w(w[1215:1184]),
        .out_w_delayed(out_w[1215:1184])
    );

    w_16_63 #(  // w38, inputs should be aligned
        .DELAY_DIST_16(21),  // w22, delay 21 cycles
        .DELAY_DIST_15(21),  // w23, delay 21 cycles
        .DELAY_DIST_7(9),  // w31, delay 9 cycles
        .DELAY_DIST_2(0),  // w36, delay 0 cycles
        .DELAY_OUT_W(116)
    ) w_38_inst( 
        .clk(clk),
        .dist_16(w[735:704]),  // w22
        .dist_15(w[767:736]),  // w23
        .dist_7(w[1023:992]),  // w31
        .dist_2(w[1183:1152]),  // w36
        .out_w(w[1247:1216]),
        .out_w_delayed(out_w[1247:1216])
    );

    w_16_63 #(  // w39, inputs should be aligned
        .DELAY_DIST_16(21),  // w23, delay 21 cycles
        .DELAY_DIST_15(18),  // w24, delay 18 cycles
        .DELAY_DIST_7(6),  // w32, delay 6 cycles
        .DELAY_DIST_2(0),  // w37, delay 0 cycles
        .DELAY_OUT_W(120)
    ) w_39_inst( 
        .clk(clk),
        .dist_16(w[767:736]),  // w23
        .dist_15(w[799:768]),  // w24
        .dist_7(w[1055:1024]),  // w32
        .dist_2(w[1215:1184]),  // w37
        .out_w(w[1279:1248]),
        .out_w_delayed(out_w[1279:1248])
    );

    w_16_63 #(  // w40, inputs should be aligned
        .DELAY_DIST_16(21),  // w24, delay 21 cycles
        .DELAY_DIST_15(21),  // w25, delay 21 cycles
        .DELAY_DIST_7(9),  // w33, delay 9 cycles
        .DELAY_DIST_2(0),  // w38, delay 0 cycles
        .DELAY_OUT_W(121)
    ) w_40_inst( 
        .clk(clk),
        .dist_16(w[799:768]),  // w24
        .dist_15(w[831:800]),  // w25
        .dist_7(w[1087:1056]),  // w33
        .dist_2(w[1247:1216]),  // w38
        .out_w(w[1311:1280]),
        .out_w_delayed(out_w[1311:1280])
    );

    w_16_63 #(  // w41, inputs should be aligned
        .DELAY_DIST_16(21),  // w25, delay 21 cycles
        .DELAY_DIST_15(18),  // w26, delay 18 cycles
        .DELAY_DIST_7(6),  // w34, delay 6 cycles
        .DELAY_DIST_2(0),  // w39, delay 0 cycles
        .DELAY_OUT_W(125)
    ) w_41_inst( 
        .clk(clk),
        .dist_16(w[831:800]),  // w25
        .dist_15(w[863:832]),  // w26
        .dist_7(w[1119:1088]),  // w34
        .dist_2(w[1279:1248]),  // w39
        .out_w(w[1343:1312]),
        .out_w_delayed(out_w[1343:1312])
    );

    w_16_63 #(  // w42, inputs should be aligned
        .DELAY_DIST_16(21),  // w26, delay 21 cycles
        .DELAY_DIST_15(21),  // w27, delay 21 cycles
        .DELAY_DIST_7(9),  // w35, delay 9 cycles
        .DELAY_DIST_2(0),  // w40, delay 0 cycles
        .DELAY_OUT_W(126)
    ) w_42_inst( 
        .clk(clk),
        .dist_16(w[863:832]),  // w26
        .dist_15(w[895:864]),  // w27
        .dist_7(w[1151:1120]),  // w35
        .dist_2(w[1311:1280]),  // w40
        .out_w(w[1375:1344]),
        .out_w_delayed(out_w[1375:1344])
    );

    w_16_63 #(  // w43, inputs should be aligned
        .DELAY_DIST_16(21),  // w27, delay 21 cycles
        .DELAY_DIST_15(18),  // w28, delay 18 cycles
        .DELAY_DIST_7(6),  // w36, delay 6 cycles
        .DELAY_DIST_2(0),  // w41, delay 0 cycles
        .DELAY_OUT_W(130)
    ) w_43_inst( 
        .clk(clk),
        .dist_16(w[895:864]),  // w27
        .dist_15(w[927:896]),  // w28
        .dist_7(w[1183:1152]),  // w36
        .dist_2(w[1343:1312]),  // w41
        .out_w(w[1407:1376]),
        .out_w_delayed(out_w[1407:1376])
    );

    w_16_63 #(  // w44, inputs should be aligned
        .DELAY_DIST_16(21),  // w28, delay 21 cycles
        .DELAY_DIST_15(21),  // w29, delay 21 cycles
        .DELAY_DIST_7(9),  // w37, delay 9 cycles
        .DELAY_DIST_2(0),  // w42, delay 0 cycles
        .DELAY_OUT_W(131)
    ) w_44_inst( 
        .clk(clk),
        .dist_16(w[927:896]),  // w28
        .dist_15(w[959:928]),  // w29
        .dist_7(w[1215:1184]),  // w37
        .dist_2(w[1375:1344]),  // w42
        .out_w(w[1439:1408]),
        .out_w_delayed(out_w[1439:1408])
    );

    w_16_63 #(  // w45, inputs should be aligned
        .DELAY_DIST_16(21),  // w29, delay 21 cycles
        .DELAY_DIST_15(18),  // w30, delay 18 cycles
        .DELAY_DIST_7(6),  // w38, delay 6 cycles
        .DELAY_DIST_2(0),  // w43, delay 0 cycles
        .DELAY_OUT_W(135)
    ) w_45_inst( 
        .clk(clk),
        .dist_16(w[959:928]),  // w29
        .dist_15(w[991:960]),  // w30
        .dist_7(w[1247:1216]),  // w38
        .dist_2(w[1407:1376]),  // w43
        .out_w(w[1471:1440]),
        .out_w_delayed(out_w[1471:1440])
    );

    w_16_63 #(  // w46, inputs should be aligned
        .DELAY_DIST_16(21),  // w30, delay 21 cycles
        .DELAY_DIST_15(21),  // w31, delay 21 cycles
        .DELAY_DIST_7(9),  // w39, delay 9 cycles
        .DELAY_DIST_2(0),  // w44, delay 0 cycles
        .DELAY_OUT_W(136)
    ) w_46_inst( 
        .clk(clk),
        .dist_16(w[991:960]),  // w30
        .dist_15(w[1023:992]),  // w31
        .dist_7(w[1279:1248]),  // w39
        .dist_2(w[1439:1408]),  // w44
        .out_w(w[1503:1472]),
        .out_w_delayed(out_w[1503:1472])
    );

    w_16_63 #(  // w47, inputs should be aligned
        .DELAY_DIST_16(21),  // w31, delay 21 cycles
        .DELAY_DIST_15(18),  // w32, delay 18 cycles
        .DELAY_DIST_7(6),  // w40, delay 6 cycles
        .DELAY_DIST_2(0),  // w45, delay 0 cycles
        .DELAY_OUT_W(140)
    ) w_47_inst( 
        .clk(clk),
        .dist_16(w[1023:992]),  // w31
        .dist_15(w[1055:1024]),  // w32
        .dist_7(w[1311:1280]),  // w40
        .dist_2(w[1471:1440]),  // w45
        .out_w(w[1535:1504]),
        .out_w_delayed(out_w[1535:1504])
    );

    w_16_63 #(  // w48, inputs should be aligned
        .DELAY_DIST_16(21),  // w32, delay 21 cycles
        .DELAY_DIST_15(21),  // w33, delay 21 cycles
        .DELAY_DIST_7(9),  // w41, delay 9 cycles
        .DELAY_DIST_2(0),  // w46, delay 0 cycles
        .DELAY_OUT_W(141)
    ) w_48_inst( 
        .clk(clk),
        .dist_16(w[1055:1024]),  // w32
        .dist_15(w[1087:1056]),  // w33
        .dist_7(w[1343:1312]),  // w41
        .dist_2(w[1503:1472]),  // w46
        .out_w(w[1567:1536]),
        .out_w_delayed(out_w[1567:1536])
    );

    w_16_63 #(  // w49, inputs should be aligned
        .DELAY_DIST_16(21),  // w33, delay 21 cycles
        .DELAY_DIST_15(18),  // w34, delay 18 cycles
        .DELAY_DIST_7(6),  // w42, delay 6 cycles
        .DELAY_DIST_2(0),  // w47, delay 0 cycles
        .DELAY_OUT_W(145)
    ) w_49_inst( 
        .clk(clk),
        .dist_16(w[1087:1056]),  // w33
        .dist_15(w[1119:1088]),  // w34
        .dist_7(w[1375:1344]),  // w42
        .dist_2(w[1535:1504]),  // w47
        .out_w(w[1599:1568]),
        .out_w_delayed(out_w[1599:1568])
    );

    w_16_63 #(  // w50, inputs should be aligned
        .DELAY_DIST_16(21),  // w34, delay 21 cycles
        .DELAY_DIST_15(21),  // w35, delay 21 cycles
        .DELAY_DIST_7(9),  // w43, delay 9 cycles
        .DELAY_DIST_2(0),  // w48, delay 0 cycles
        .DELAY_OUT_W(146)
    ) w_50_inst( 
        .clk(clk),
        .dist_16(w[1119:1088]),  // w34
        .dist_15(w[1151:1120]),  // w35
        .dist_7(w[1407:1376]),  // w43
        .dist_2(w[1567:1536]),  // w48
        .out_w(w[1631:1600]),
        .out_w_delayed(out_w[1631:1600])
    );

    w_16_63 #(  // w51, inputs should be aligned
        .DELAY_DIST_16(21),  // w35, delay 21 cycles
        .DELAY_DIST_15(18),  // w36, delay 18 cycles
        .DELAY_DIST_7(6),  // w44, delay 6 cycles
        .DELAY_DIST_2(0),  // w49, delay 0 cycles
        .DELAY_OUT_W(150)
    ) w_51_inst( 
        .clk(clk),
        .dist_16(w[1151:1120]),  // w35
        .dist_15(w[1183:1152]),  // w36
        .dist_7(w[1439:1408]),  // w44
        .dist_2(w[1599:1568]),  // w49
        .out_w(w[1663:1632]),
        .out_w_delayed(out_w[1663:1632])
    );

    w_16_63 #(  // w52, inputs should be aligned
        .DELAY_DIST_16(21),  // w36, delay 21 cycles
        .DELAY_DIST_15(21),  // w37, delay 21 cycles
        .DELAY_DIST_7(9),  // w45, delay 9 cycles
        .DELAY_DIST_2(0),  // w50, delay 0 cycles
        .DELAY_OUT_W(151)
    ) w_52_inst( 
        .clk(clk),
        .dist_16(w[1183:1152]),  // w36
        .dist_15(w[1215:1184]),  // w37
        .dist_7(w[1471:1440]),  // w45
        .dist_2(w[1631:1600]),  // w50
        .out_w(w[1695:1664]),
        .out_w_delayed(out_w[1695:1664])
    );

    w_16_63 #(  // w53, inputs should be aligned
        .DELAY_DIST_16(21),  // w37, delay 21 cycles
        .DELAY_DIST_15(18),  // w38, delay 18 cycles
        .DELAY_DIST_7(6),  // w46, delay 6 cycles
        .DELAY_DIST_2(0),  // w51, delay 0 cycles
        .DELAY_OUT_W(155)
    ) w_53_inst( 
        .clk(clk),
        .dist_16(w[1215:1184]),  // w37
        .dist_15(w[1247:1216]),  // w38
        .dist_7(w[1503:1472]),  // w46
        .dist_2(w[1663:1632]),  // w51
        .out_w(w[1727:1696]),
        .out_w_delayed(out_w[1727:1696])
    );

    w_16_63 #(  // w54, inputs should be aligned
        .DELAY_DIST_16(21),  // w38, delay 21 cycles
        .DELAY_DIST_15(21),  // w39, delay 21 cycles
        .DELAY_DIST_7(9),  // w47, delay 9 cycles
        .DELAY_DIST_2(0),  // w52, delay 0 cycles
        .DELAY_OUT_W(156)
    ) w_54_inst( 
        .clk(clk),
        .dist_16(w[1247:1216]),  // w38
        .dist_15(w[1279:1248]),  // w39
        .dist_7(w[1535:1504]),  // w47
        .dist_2(w[1695:1664]),  // w52
        .out_w(w[1759:1728]),
        .out_w_delayed(out_w[1759:1728])
    );

    w_16_63 #(  // w55, inputs should be aligned
        .DELAY_DIST_16(21),  // w39, delay 21 cycles
        .DELAY_DIST_15(18),  // w40, delay 18 cycles
        .DELAY_DIST_7(6),  // w48, delay 6 cycles
        .DELAY_DIST_2(0),  // w53, delay 0 cycles
        .DELAY_OUT_W(160)
    ) w_55_inst( 
        .clk(clk),
        .dist_16(w[1279:1248]),  // w39
        .dist_15(w[1311:1280]),  // w40
        .dist_7(w[1567:1536]),  // w48
        .dist_2(w[1727:1696]),  // w53
        .out_w(w[1791:1760]),
        .out_w_delayed(out_w[1791:1760])
    );

    w_16_63 #(  // w56, inputs should be aligned
        .DELAY_DIST_16(21),  // w40, delay 21 cycles
        .DELAY_DIST_15(21),  // w41, delay 21 cycles
        .DELAY_DIST_7(9),  // w49, delay 9 cycles
        .DELAY_DIST_2(0),  // w54, delay 0 cycles
        .DELAY_OUT_W(161)
    ) w_56_inst( 
        .clk(clk),
        .dist_16(w[1311:1280]),  // w40
        .dist_15(w[1343:1312]),  // w41
        .dist_7(w[1599:1568]),  // w49
        .dist_2(w[1759:1728]),  // w54
        .out_w(w[1823:1792]),
        .out_w_delayed(out_w[1823:1792])
    );

    w_16_63 #(  // w57, inputs should be aligned
        .DELAY_DIST_16(21),  // w41, delay 21 cycles
        .DELAY_DIST_15(18),  // w42, delay 18 cycles
        .DELAY_DIST_7(6),  // w50, delay 6 cycles
        .DELAY_DIST_2(0),  // w55, delay 0 cycles
        .DELAY_OUT_W(165)
    ) w_57_inst( 
        .clk(clk),
        .dist_16(w[1343:1312]),  // w41
        .dist_15(w[1375:1344]),  // w42
        .dist_7(w[1631:1600]),  // w50
        .dist_2(w[1791:1760]),  // w55
        .out_w(w[1855:1824]),
        .out_w_delayed(out_w[1855:1824])
    );

    w_16_63 #(  // w58, inputs should be aligned
        .DELAY_DIST_16(21),  // w42, delay 21 cycles
        .DELAY_DIST_15(21),  // w43, delay 21 cycles
        .DELAY_DIST_7(9),  // w51, delay 9 cycles
        .DELAY_DIST_2(0),  // w56, delay 0 cycles
        .DELAY_OUT_W(166)
    ) w_58_inst( 
        .clk(clk),
        .dist_16(w[1375:1344]),  // w42
        .dist_15(w[1407:1376]),  // w43
        .dist_7(w[1663:1632]),  // w51
        .dist_2(w[1823:1792]),  // w56
        .out_w(w[1887:1856]),
        .out_w_delayed(out_w[1887:1856])
    );

    w_16_63 #(  // w59, inputs should be aligned
        .DELAY_DIST_16(21),  // w43, delay 21 cycles
        .DELAY_DIST_15(18),  // w44, delay 18 cycles
        .DELAY_DIST_7(6),  // w52, delay 6 cycles
        .DELAY_DIST_2(0),  // w57, delay 0 cycles
        .DELAY_OUT_W(170)
    ) w_59_inst( 
        .clk(clk),
        .dist_16(w[1407:1376]),  // w43
        .dist_15(w[1439:1408]),  // w44
        .dist_7(w[1695:1664]),  // w52
        .dist_2(w[1855:1824]),  // w57
        .out_w(w[1919:1888]),
        .out_w_delayed(out_w[1919:1888])
    );

    w_16_63 #(  // w60, inputs should be aligned
        .DELAY_DIST_16(21),  // w44, delay 21 cycles
        .DELAY_DIST_15(21),  // w45, delay 21 cycles
        .DELAY_DIST_7(9),  // w53, delay 9 cycles
        .DELAY_DIST_2(0),  // w58, delay 0 cycles
        .DELAY_OUT_W(171)
    ) w_60_inst( 
        .clk(clk),
        .dist_16(w[1439:1408]),  // w44
        .dist_15(w[1471:1440]),  // w45
        .dist_7(w[1727:1696]),  // w53
        .dist_2(w[1887:1856]),  // w58
        .out_w(w[1951:1920]),
        .out_w_delayed(out_w[1951:1920])
    );

    w_16_63 #(  // w61, inputs should be aligned
        .DELAY_DIST_16(21),  // w45, delay 21 cycles
        .DELAY_DIST_15(18),  // w46, delay 18 cycles
        .DELAY_DIST_7(6),  // w54, delay 6 cycles
        .DELAY_DIST_2(0),  // w59, delay 0 cycles
        .DELAY_OUT_W(175)
    ) w_61_inst( 
        .clk(clk),
        .dist_16(w[1471:1440]),  // w45
        .dist_15(w[1503:1472]),  // w46
        .dist_7(w[1759:1728]),  // w54
        .dist_2(w[1919:1888]),  // w59
        .out_w(w[1983:1952]),
        .out_w_delayed(out_w[1983:1952])
    );

    w_16_63 #(  // w62, inputs should be aligned
        .DELAY_DIST_16(21),  // w46, delay 21 cycles
        .DELAY_DIST_15(21),  // w47, delay 21 cycles
        .DELAY_DIST_7(9),  // w55, delay 9 cycles
        .DELAY_DIST_2(0),  // w60, delay 0 cycles
        .DELAY_OUT_W(176)
    ) w_62_inst( 
        .clk(clk),
        .dist_16(w[1503:1472]),  // w46
        .dist_15(w[1535:1504]),  // w47
        .dist_7(w[1791:1760]),  // w55
        .dist_2(w[1951:1920]),  // w60
        .out_w(w[2015:1984]),
        .out_w_delayed(out_w[2015:1984])
    );

    w_16_63 #(  // w63, inputs should be aligned
        .DELAY_DIST_16(21),  // w47, delay 21 cycles
        .DELAY_DIST_15(18),  // w48, delay 18 cycles
        .DELAY_DIST_7(6),  // w56, delay 6 cycles
        .DELAY_DIST_2(0),  // w61, delay 0 cycles
        .DELAY_OUT_W(180)
    ) w_63_inst( 
        .clk(clk),
        .dist_16(w[1535:1504]),  // w47
        .dist_15(w[1567:1536]),  // w48
        .dist_7(w[1823:1792]),  // w56
        .dist_2(w[1983:1952]),  // w61
        .out_w(w[2047:2016]),
        .out_w_delayed(out_w[2047:2016])
    );

endmodule

//
// w[0..15]
//
module w_0_15 #(
    parameter DELAY_OUT_W = 0
)(
    input clk,
    input [31:0] chunk,
    output reg [31:0] out_w = 0,
    output [31:0] out_w_delayed
);
    always @(posedge clk) begin
        out_w[7:0] <= chunk[31:24];
        out_w[15:8] <= chunk[23:16];
        out_w[23:16] <= chunk[15:8];
        out_w[31:24] <= chunk[7:0];
    end

    shift_reg #(
        .DELAY(DELAY_OUT_W),
        .DATA_WIDTH(32)
    ) shift_reg_out_w(
    	.clk(clk),
        .i(out_w),
        .o(out_w_delayed)
    );
endmodule

//
// w[16..63]
//
module w_16_63 #(
    parameter DELAY_DIST_16 = 0,  // input delay of dist_16
    parameter DELAY_DIST_15 = 0,  // input delay of dist_15
    parameter DELAY_DIST_7 = 0,  // input delay of dist_7
    parameter DELAY_DIST_2 = 0,  // input delay of dist_2
    parameter DELAY_OUT_W = 0  // output delay 
)(
    input clk,
    input [31:0] dist_16,
    input [31:0] dist_15,
    input [31:0] dist_7,
    input [31:0] dist_2,
    output [31:0] out_w,
    output [31:0] out_w_delayed
);
    //
    // delayed inputs
    //
    wire [31:0] delayed_dist_16;
    wire [31:0] delayed_dist_15;
    wire [31:0] delayed_dist_7;
    wire [31:0] delayed_dist_2;

    shift_reg #(
        .DELAY(DELAY_DIST_16),
        .DATA_WIDTH(32)
    ) shift_reg_dist_16(
    	.clk(clk),
        .i(dist_16),
        .o(delayed_dist_16)
    );

    shift_reg #(
        .DELAY(DELAY_DIST_15),
        .DATA_WIDTH(32)
    ) shift_reg_dist_15(
    	.clk(clk),
        .i(dist_15),
        .o(delayed_dist_15)
    );

    shift_reg #(
        .DELAY(DELAY_DIST_7),
        .DATA_WIDTH(32)
    ) shift_reg_dist_7(
    	.clk(clk),
        .i(dist_7),
        .o(delayed_dist_7)
    );

    shift_reg #(
        .DELAY(DELAY_DIST_2),
        .DATA_WIDTH(32)
    ) shift_reg_dist_2(
    	.clk(clk),
        .i(dist_2),
        .o(delayed_dist_2)
    );

    //
    // Pipeline stages
    //
    // stage1. s0, s1
    reg [31:0] s1_s0 = 0;
    reg [31:0] s1_s1 = 0;
    reg [31:0] s1_dist_16 = 0;
    reg [31:0] s1_dist_7 = 0;

    always @(posedge clk) begin
        s1_s0 <= {delayed_dist_15[6:0], delayed_dist_15[31:7]} ^ {delayed_dist_15[17:0], delayed_dist_15[31:18]} ^ {{3{1'b0}}, delayed_dist_15[31:3]};
        s1_s1 <= {delayed_dist_2[16:0], delayed_dist_2[31:17]} ^ {delayed_dist_2[18:0], delayed_dist_2[31:19]} ^ {{10{1'b0}}, delayed_dist_2[31:10]};
        s1_dist_16 <= delayed_dist_16;
        s1_dist_7 <= delayed_dist_7;
    end

    // stage2. sum_s, sum_w
    reg [31:0] s2_sum_s = 0;
    reg [31:0] s2_sum_w = 0;

    always @(posedge clk) begin
        s2_sum_s <= s1_s0+s1_s1;
        s2_sum_w <= s1_dist_16+s1_dist_7;
    end

    // stage3. w
    reg [31:0] s3_out_w = 0;

    always @(posedge clk) begin
        s3_out_w <= s2_sum_s+s2_sum_w;
    end

    assign out_w = s3_out_w;

    //
    // delayed output
    //
    shift_reg #(
        .DELAY(DELAY_OUT_W),
        .DATA_WIDTH(32)
    ) shift_reg_out_w(
    	.clk(clk),
        .i(s3_out_w),
        .o(out_w_delayed)
    );
endmodule
